library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity program_counter is
    port(
        clk : in std_logic;
        rst : in std_logic
    );
end entity program_counter;

architecture RTL of program_counter is
    
begin

end architecture RTL;
